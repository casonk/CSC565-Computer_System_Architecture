
module bit_memory_unit_test;

	// Inputs
	reg inbit_0;
	// reg inbit_1;
	reg load_flag;

	// Outputs
	wire outbit_0;
	// wire carry_out; 
	// wire borrow_out;

	// Instantiate the Unit Under Test (UUT)
	bit_memory_unit uut (
		.inbit_0(inbit_0), 
		// .inbit_1(inbit_1),
		.load_flag (load_flag),
		.outbit_0(outbit_0)
		// .carry_out(carry_out)
		// .borrow_out(borrow_out)
		
	);

	initial begin
		// Initialize Inputs
		inbit_0 = 0;
		// inbit_1 = 0;
		load_flag = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here: 100 INPUTS

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 0;
        #100;
        

        inbit_0 = 0;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

        inbit_0 = 1;
        // inbit_1 = ;
		load_flag = 1;
        #100;
        

    end
endmodule
