
module module_test;

	// Inputs
	reg inx;
	reg iny;

	// Outputs
	wire ouz;

	// Instantiate the Unit Under Test (UUT)
	module uut (
		.inx(inx), 
		.iny(iny), 
		.ouz(ouz)
	);

	initial begin
		// Initialize Inputs
		inx = 00000000;
		iny = 00000000;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here: 1000 INPUTS

        inx = 01011000;
        iny = 01000110;
        #100;


        inx = 00011101;
        iny = 11111111;
        #100;


        inx = 11101101;
        iny = 11110100;
        #100;


        inx = 00000000;
        iny = 10010010;
        #100;


        inx = 10000001;
        iny = 01100101;
        #100;


        inx = 01000111;
        iny = 11011111;
        #100;


        inx = 10100100;
        iny = 10001001;
        #100;


        inx = 00010111;
        iny = 11010110;
        #100;


        inx = 11010100;
        iny = 10001101;
        #100;


        inx = 00010010;
        iny = 00001101;
        #100;


        inx = 00001010;
        iny = 00000010;
        #100;


        inx = 01011100;
        iny = 00001110;
        #100;


        inx = 00000110;
        iny = 01111001;
        #100;


        inx = 01110011;
        iny = 11100000;
        #100;


        inx = 10110010;
        iny = 11000010;
        #100;


        inx = 10001100;
        iny = 11100010;
        #100;


        inx = 00101111;
        iny = 10110101;
        #100;


        inx = 10110101;
        iny = 11000010;
        #100;


        inx = 01110110;
        iny = 11010111;
        #100;


        inx = 11111101;
        iny = 00011000;
        #100;


        inx = 01011110;
        iny = 11011000;
        #100;


        inx = 01011111;
        iny = 01111111;
        #100;


        inx = 01010111;
        iny = 11101111;
        #100;


        inx = 10000010;
        iny = 10110011;
        #100;


        inx = 01101000;
        iny = 00111011;
        #100;


        inx = 00101000;
        iny = 00000110;
        #100;


        inx = 10101101;
        iny = 11101111;
        #100;


        inx = 11001101;
        iny = 01111110;
        #100;


        inx = 11101011;
        iny = 10110011;
        #100;


        inx = 10011111;
        iny = 10100101;
        #100;


        inx = 01001000;
        iny = 01100011;
        #100;


        inx = 00000000;
        iny = 11110010;
        #100;


        inx = 01000110;
        iny = 01110111;
        #100;


        inx = 11110111;
        iny = 10110011;
        #100;


        inx = 11111001;
        iny = 01101000;
        #100;


        inx = 00001101;
        iny = 10111010;
        #100;


        inx = 00101001;
        iny = 11101100;
        #100;


        inx = 11110101;
        iny = 01100100;
        #100;


        inx = 00001011;
        iny = 10010101;
        #100;


        inx = 11111010;
        iny = 10110110;
        #100;


        inx = 01010011;
        iny = 10001010;
        #100;


        inx = 00010110;
        iny = 11001001;
        #100;


        inx = 01111000;
        iny = 11000101;
        #100;


        inx = 00101100;
        iny = 00110100;
        #100;


        inx = 01010011;
        iny = 00010001;
        #100;


        inx = 00001000;
        iny = 00000101;
        #100;


        inx = 10001100;
        iny = 01101100;
        #100;


        inx = 01110111;
        iny = 00001100;
        #100;


        inx = 00100101;
        iny = 01111000;
        #100;


        inx = 11010011;
        iny = 10001111;
        #100;


        inx = 11110001;
        iny = 10010010;
        #100;


        inx = 11001111;
        iny = 11001111;
        #100;


        inx = 11001010;
        iny = 10101001;
        #100;


        inx = 11011010;
        iny = 00111101;
        #100;


        inx = 00101111;
        iny = 01100111;
        #100;


        inx = 11011111;
        iny = 01001100;
        #100;


        inx = 11110000;
        iny = 10001111;
        #100;


        inx = 10011010;
        iny = 11010010;
        #100;


        inx = 01001011;
        iny = 11000110;
        #100;


        inx = 11010010;
        iny = 01110001;
        #100;


        inx = 00001101;
        iny = 10000111;
        #100;


        inx = 01011011;
        iny = 01111101;
        #100;


        inx = 00100000;
        iny = 00100100;
        #100;


        inx = 11111111;
        iny = 10010011;
        #100;


        inx = 00110010;
        iny = 11100101;
        #100;


        inx = 11111110;
        iny = 11111100;
        #100;


        inx = 00110010;
        iny = 10011001;
        #100;


        inx = 11110011;
        iny = 11000100;
        #100;


        inx = 00000100;
        iny = 01100000;
        #100;


        inx = 00011010;
        iny = 10010011;
        #100;


        inx = 00101001;
        iny = 00010111;
        #100;


        inx = 10000001;
        iny = 01111110;
        #100;


        inx = 10111100;
        iny = 01101100;
        #100;


        inx = 01110110;
        iny = 00010100;
        #100;


        inx = 00011011;
        iny = 11101000;
        #100;


        inx = 00101100;
        iny = 10001010;
        #100;


        inx = 10111001;
        iny = 01100010;
        #100;


        inx = 10111100;
        iny = 01111111;
        #100;


        inx = 11011101;
        iny = 10001101;
        #100;


        inx = 01101101;
        iny = 00111000;
        #100;


        inx = 10010010;
        iny = 00010111;
        #100;


        inx = 00110000;
        iny = 00011111;
        #100;


        inx = 00110011;
        iny = 01110010;
        #100;


        inx = 00000001;
        iny = 11010010;
        #100;


        inx = 00100100;
        iny = 01111011;
        #100;


        inx = 11111111;
        iny = 10101111;
        #100;


        inx = 10111000;
        iny = 10010011;
        #100;


        inx = 11110010;
        iny = 00010100;
        #100;


        inx = 11100001;
        iny = 10101000;
        #100;


        inx = 11001000;
        iny = 11000000;
        #100;


        inx = 00011010;
        iny = 00001000;
        #100;


        inx = 01100011;
        iny = 00110011;
        #100;


        inx = 11100000;
        iny = 11110000;
        #100;


        inx = 00000110;
        iny = 11000100;
        #100;


        inx = 00010010;
        iny = 01011111;
        #100;


        inx = 11101100;
        iny = 11101011;
        #100;


        inx = 00110111;
        iny = 11011100;
        #100;


        inx = 10000111;
        iny = 01010100;
        #100;


        inx = 10110000;
        iny = 00000001;
        #100;


        inx = 11110101;
        iny = 00011100;
        #100;


        inx = 00101111;
        iny = 00101010;
        #100;


        inx = 11100101;
        iny = 10101001;
        #100;


        inx = 11100110;
        iny = 00111110;
        #100;


        inx = 00011100;
        iny = 11100101;
        #100;


        inx = 11011000;
        iny = 10010010;
        #100;


        inx = 11100001;
        iny = 00100000;
        #100;


        inx = 10001000;
        iny = 10110001;
        #100;


        inx = 10110100;
        iny = 10010101;
        #100;


        inx = 00001011;
        iny = 11110100;
        #100;


        inx = 10011110;
        iny = 11000011;
        #100;


        inx = 01001101;
        iny = 01000010;
        #100;


        inx = 10101011;
        iny = 01111010;
        #100;


        inx = 11001010;
        iny = 11010010;
        #100;


        inx = 11000010;
        iny = 11000100;
        #100;


        inx = 11111000;
        iny = 00011000;
        #100;


        inx = 10111001;
        iny = 10111010;
        #100;


        inx = 10001110;
        iny = 00011111;
        #100;


        inx = 00011111;
        iny = 11001001;
        #100;


        inx = 10000100;
        iny = 00100011;
        #100;


        inx = 00110011;
        iny = 10011100;
        #100;


        inx = 11000001;
        iny = 01110010;
        #100;


        inx = 10000110;
        iny = 00100101;
        #100;


        inx = 01011010;
        iny = 01101011;
        #100;


        inx = 00000100;
        iny = 10011000;
        #100;


        inx = 01000110;
        iny = 10010110;
        #100;


        inx = 00011011;
        iny = 00110011;
        #100;


        inx = 00011011;
        iny = 10110110;
        #100;


        inx = 01111101;
        iny = 10110011;
        #100;


        inx = 00000010;
        iny = 10111111;
        #100;


        inx = 01000011;
        iny = 00000110;
        #100;


        inx = 01100010;
        iny = 11001011;
        #100;


        inx = 10000100;
        iny = 10101011;
        #100;


        inx = 00110000;
        iny = 00110110;
        #100;


        inx = 01010001;
        iny = 00011101;
        #100;


        inx = 11010010;
        iny = 10110101;
        #100;


        inx = 01011110;
        iny = 10000011;
        #100;


        inx = 00001000;
        iny = 10110110;
        #100;


        inx = 01011000;
        iny = 11100001;
        #100;


        inx = 11010111;
        iny = 11101000;
        #100;


        inx = 11111101;
        iny = 11011000;
        #100;


        inx = 11001100;
        iny = 01000001;
        #100;


        inx = 11110101;
        iny = 11100110;
        #100;


        inx = 11101001;
        iny = 01110010;
        #100;


        inx = 00110111;
        iny = 00011011;
        #100;


        inx = 10110011;
        iny = 00101011;
        #100;


        inx = 11101101;
        iny = 11101111;
        #100;


        inx = 10000011;
        iny = 10100010;
        #100;


        inx = 11111000;
        iny = 11010100;
        #100;


        inx = 11011000;
        iny = 00010001;
        #100;


        inx = 00100000;
        iny = 01100110;
        #100;


        inx = 11010110;
        iny = 11001010;
        #100;


        inx = 00111110;
        iny = 10110110;
        #100;


        inx = 11001001;
        iny = 11100001;
        #100;


        inx = 01010110;
        iny = 01000101;
        #100;


        inx = 01100101;
        iny = 01010000;
        #100;


        inx = 00001110;
        iny = 01001100;
        #100;


        inx = 00110111;
        iny = 00010101;
        #100;


        inx = 10111110;
        iny = 00010001;
        #100;


        inx = 11001110;
        iny = 00111110;
        #100;


        inx = 00000111;
        iny = 01111000;
        #100;


        inx = 01110110;
        iny = 01101001;
        #100;


        inx = 10111000;
        iny = 10001000;
        #100;


        inx = 00110100;
        iny = 00111100;
        #100;


        inx = 11001011;
        iny = 00000001;
        #100;


        inx = 11101011;
        iny = 00011101;
        #100;


        inx = 11111101;
        iny = 11001010;
        #100;


        inx = 11001110;
        iny = 01001111;
        #100;


        inx = 00111001;
        iny = 10110110;
        #100;


        inx = 01111110;
        iny = 11111011;
        #100;


        inx = 10010110;
        iny = 10100111;
        #100;


        inx = 10100100;
        iny = 01010111;
        #100;


        inx = 00110001;
        iny = 10000001;
        #100;


        inx = 10101010;
        iny = 11010101;
        #100;


        inx = 01000100;
        iny = 00101110;
        #100;


        inx = 10000111;
        iny = 00110100;
        #100;


        inx = 01110001;
        iny = 10111101;
        #100;


        inx = 00001000;
        iny = 10110111;
        #100;


        inx = 01011100;
        iny = 11011011;
        #100;


        inx = 10011011;
        iny = 00010001;
        #100;


        inx = 10001011;
        iny = 01010100;
        #100;


        inx = 01010010;
        iny = 10110111;
        #100;


        inx = 01111000;
        iny = 10010100;
        #100;


        inx = 11010010;
        iny = 10100001;
        #100;


        inx = 01101000;
        iny = 10010000;
        #100;


        inx = 11110101;
        iny = 10001110;
        #100;


        inx = 10010010;
        iny = 10010100;
        #100;


        inx = 10110101;
        iny = 11011011;
        #100;


        inx = 00110000;
        iny = 00001100;
        #100;


        inx = 10101011;
        iny = 10010100;
        #100;


        inx = 01101010;
        iny = 11001010;
        #100;


        inx = 01010001;
        iny = 01110110;
        #100;


        inx = 00100100;
        iny = 11010101;
        #100;


        inx = 01000101;
        iny = 10011100;
        #100;


        inx = 01011000;
        iny = 11011010;
        #100;


        inx = 00001000;
        iny = 01110000;
        #100;


        inx = 10110111;
        iny = 00011010;
        #100;


        inx = 11000001;
        iny = 10100011;
        #100;


        inx = 11000010;
        iny = 01110010;
        #100;


        inx = 11110111;
        iny = 00000100;
        #100;


        inx = 00011011;
        iny = 10011010;
        #100;


        inx = 01111000;
        iny = 00100000;
        #100;


        inx = 00101111;
        iny = 00000100;
        #100;


        inx = 10100011;
        iny = 01101011;
        #100;


        inx = 01001011;
        iny = 01100001;
        #100;


        inx = 11011011;
        iny = 10011001;
        #100;


        inx = 10111101;
        iny = 11110111;
        #100;


        inx = 00000101;
        iny = 11010011;
        #100;


        inx = 01110011;
        iny = 01001101;
        #100;


        inx = 11111111;
        iny = 01011001;
        #100;


        inx = 01011100;
        iny = 10100010;
        #100;


        inx = 01111001;
        iny = 11110100;
        #100;


        inx = 10000110;
        iny = 11100001;
        #100;


        inx = 00010010;
        iny = 11011000;
        #100;


        inx = 01000001;
        iny = 10001010;
        #100;


        inx = 10001101;
        iny = 11001101;
        #100;


        inx = 01010001;
        iny = 10011011;
        #100;


        inx = 01111000;
        iny = 00011000;
        #100;


        inx = 10101110;
        iny = 01010111;
        #100;


        inx = 00101011;
        iny = 11010000;
        #100;


        inx = 00110011;
        iny = 10001010;
        #100;


        inx = 11011011;
        iny = 11100001;
        #100;


        inx = 01111110;
        iny = 11001100;
        #100;


        inx = 11110111;
        iny = 00110100;
        #100;


        inx = 11011100;
        iny = 11010100;
        #100;


        inx = 11111010;
        iny = 00001110;
        #100;


        inx = 11101100;
        iny = 00101100;
        #100;


        inx = 01010100;
        iny = 10101010;
        #100;


        inx = 11010000;
        iny = 00000100;
        #100;


        inx = 00101100;
        iny = 10001010;
        #100;


        inx = 10100011;
        iny = 10100011;
        #100;


        inx = 00000010;
        iny = 01110010;
        #100;


        inx = 01100101;
        iny = 10001100;
        #100;


        inx = 00010110;
        iny = 11011110;
        #100;


        inx = 11110110;
        iny = 11011110;
        #100;


        inx = 10101011;
        iny = 00011100;
        #100;


        inx = 01010010;
        iny = 00001000;
        #100;


        inx = 11101100;
        iny = 00110000;
        #100;


        inx = 00000110;
        iny = 11100101;
        #100;


        inx = 10100110;
        iny = 11110001;
        #100;


        inx = 10000100;
        iny = 11101101;
        #100;


        inx = 01011010;
        iny = 01100011;
        #100;


        inx = 10101001;
        iny = 01010110;
        #100;


        inx = 01001000;
        iny = 10010011;
        #100;


        inx = 00001010;
        iny = 11000011;
        #100;


        inx = 10000100;
        iny = 01010010;
        #100;


        inx = 00111101;
        iny = 01001000;
        #100;


        inx = 11000111;
        iny = 10001110;
        #100;


        inx = 01010100;
        iny = 01110000;
        #100;


        inx = 01000111;
        iny = 11110011;
        #100;


        inx = 10101100;
        iny = 01111001;
        #100;


        inx = 11000001;
        iny = 10011000;
        #100;


        inx = 10110110;
        iny = 01100100;
        #100;


        inx = 00101100;
        iny = 00111110;
        #100;


        inx = 01010010;
        iny = 11110000;
        #100;


        inx = 10100000;
        iny = 00110101;
        #100;


        inx = 10111010;
        iny = 00011000;
        #100;


        inx = 11011000;
        iny = 11111100;
        #100;


        inx = 00010000;
        iny = 10000010;
        #100;


        inx = 00011011;
        iny = 11010101;
        #100;


        inx = 01010010;
        iny = 10100001;
        #100;


        inx = 11011111;
        iny = 01100010;
        #100;


        inx = 11000111;
        iny = 10010110;
        #100;


        inx = 01101100;
        iny = 01011011;
        #100;


        inx = 10001111;
        iny = 00010010;
        #100;


        inx = 01111000;
        iny = 11111111;
        #100;


        inx = 11001011;
        iny = 11110111;
        #100;


        inx = 01001111;
        iny = 11100101;
        #100;


        inx = 01100011;
        iny = 00110011;
        #100;


        inx = 00011011;
        iny = 00110010;
        #100;


        inx = 01001000;
        iny = 11010000;
        #100;


        inx = 11110101;
        iny = 11100110;
        #100;


        inx = 11101011;
        iny = 01100100;
        #100;


        inx = 11000011;
        iny = 11011010;
        #100;


        inx = 11010100;
        iny = 11101010;
        #100;


        inx = 01001110;
        iny = 11100110;
        #100;


        inx = 10110001;
        iny = 11100101;
        #100;


        inx = 01110111;
        iny = 11100010;
        #100;


        inx = 11000110;
        iny = 11010101;
        #100;


        inx = 10001010;
        iny = 10001010;
        #100;


        inx = 00000000;
        iny = 11110101;
        #100;


        inx = 10011111;
        iny = 10010011;
        #100;


        inx = 01100000;
        iny = 11000101;
        #100;


        inx = 01101010;
        iny = 00100110;
        #100;


        inx = 11011110;
        iny = 11000100;
        #100;


        inx = 11000111;
        iny = 00010110;
        #100;


        inx = 10011000;
        iny = 11000110;
        #100;


        inx = 10000011;
        iny = 11001111;
        #100;


        inx = 00101000;
        iny = 10000001;
        #100;


        inx = 00001000;
        iny = 00000101;
        #100;


        inx = 01010111;
        iny = 01101111;
        #100;


        inx = 10000111;
        iny = 01110110;
        #100;


        inx = 00101011;
        iny = 10110011;
        #100;


        inx = 00001011;
        iny = 11000001;
        #100;


        inx = 01011111;
        iny = 11100111;
        #100;


        inx = 00101001;
        iny = 01101110;
        #100;


        inx = 10101000;
        iny = 11100100;
        #100;


        inx = 10010110;
        iny = 00011000;
        #100;


        inx = 01010000;
        iny = 11000111;
        #100;


        inx = 11000001;
        iny = 00110100;
        #100;


        inx = 11101100;
        iny = 00101011;
        #100;


        inx = 01011101;
        iny = 10010010;
        #100;


        inx = 01100101;
        iny = 01110011;
        #100;


        inx = 10011111;
        iny = 01000000;
        #100;


        inx = 10011100;
        iny = 10100110;
        #100;


        inx = 10001001;
        iny = 01110110;
        #100;


        inx = 11010011;
        iny = 00010011;
        #100;


        inx = 01011011;
        iny = 11110011;
        #100;


        inx = 11001100;
        iny = 10010011;
        #100;


        inx = 00010101;
        iny = 10001110;
        #100;


        inx = 00010100;
        iny = 01110010;
        #100;


        inx = 11111011;
        iny = 00111000;
        #100;


        inx = 01101111;
        iny = 10101011;
        #100;


        inx = 11100111;
        iny = 00010000;
        #100;


        inx = 10100000;
        iny = 10010001;
        #100;


        inx = 00111110;
        iny = 00100001;
        #100;


        inx = 10100111;
        iny = 00000111;
        #100;


        inx = 01001011;
        iny = 01011010;
        #100;


        inx = 11111000;
        iny = 01011100;
        #100;


        inx = 10111011;
        iny = 00001011;
        #100;


        inx = 01101011;
        iny = 11011110;
        #100;


        inx = 01000111;
        iny = 01110001;
        #100;


        inx = 00100110;
        iny = 01001010;
        #100;


        inx = 10110000;
        iny = 01111010;
        #100;


        inx = 00101111;
        iny = 00011010;
        #100;


        inx = 10101010;
        iny = 10111101;
        #100;


        inx = 10110010;
        iny = 01010110;
        #100;


        inx = 00100111;
        iny = 11010100;
        #100;


        inx = 10101111;
        iny = 10000101;
        #100;


        inx = 01001001;
        iny = 01010011;
        #100;


        inx = 00000101;
        iny = 00100101;
        #100;


        inx = 01100101;
        iny = 01101011;
        #100;


        inx = 01110110;
        iny = 10111010;
        #100;


        inx = 11001011;
        iny = 01001100;
        #100;


        inx = 00010100;
        iny = 11111010;
        #100;


        inx = 11000000;
        iny = 11010101;
        #100;


        inx = 00111100;
        iny = 00000001;
        #100;


        inx = 10001100;
        iny = 10110010;
        #100;


        inx = 10001010;
        iny = 10100001;
        #100;


        inx = 11100001;
        iny = 00101010;
        #100;


        inx = 01111100;
        iny = 01111110;
        #100;


        inx = 01101110;
        iny = 11010101;
        #100;


        inx = 11100111;
        iny = 00001010;
        #100;


        inx = 10011101;
        iny = 01000100;
        #100;


        inx = 10110110;
        iny = 00010100;
        #100;


        inx = 01011000;
        iny = 11111101;
        #100;


        inx = 00000110;
        iny = 01001000;
        #100;


        inx = 00010111;
        iny = 00101000;
        #100;


        inx = 00000110;
        iny = 11011111;
        #100;


        inx = 00000000;
        iny = 00010100;
        #100;


        inx = 10011111;
        iny = 10000000;
        #100;


        inx = 00011111;
        iny = 11010000;
        #100;


        inx = 11001010;
        iny = 01010011;
        #100;


        inx = 01000000;
        iny = 00110010;
        #100;


        inx = 10111111;
        iny = 00110010;
        #100;


        inx = 10100011;
        iny = 01001111;
        #100;


        inx = 00111010;
        iny = 00000101;
        #100;


        inx = 10011011;
        iny = 11101110;
        #100;


        inx = 01111011;
        iny = 01010100;
        #100;


        inx = 00000000;
        iny = 10100101;
        #100;


        inx = 00010011;
        iny = 01011101;
        #100;


        inx = 01010010;
        iny = 00101010;
        #100;


        inx = 00110001;
        iny = 10011010;
        #100;


        inx = 10100101;
        iny = 00110101;
        #100;


        inx = 10000000;
        iny = 11111011;
        #100;


        inx = 00010001;
        iny = 10101101;
        #100;


        inx = 11101010;
        iny = 10010100;
        #100;


        inx = 00110100;
        iny = 00100111;
        #100;


        inx = 11011011;
        iny = 10011100;
        #100;


        inx = 01001011;
        iny = 01001100;
        #100;


        inx = 01111001;
        iny = 10000001;
        #100;


        inx = 00010111;
        iny = 10011110;
        #100;


        inx = 00100101;
        iny = 10110011;
        #100;


        inx = 00110010;
        iny = 00101110;
        #100;


        inx = 10010000;
        iny = 00011010;
        #100;


        inx = 00100001;
        iny = 01100000;
        #100;


        inx = 01011110;
        iny = 00111010;
        #100;


        inx = 10101000;
        iny = 00101010;
        #100;


        inx = 01110100;
        iny = 01110101;
        #100;


        inx = 01011101;
        iny = 10100101;
        #100;


        inx = 00010000;
        iny = 10111101;
        #100;


        inx = 10011011;
        iny = 01001111;
        #100;


        inx = 11000010;
        iny = 10000000;
        #100;


        inx = 11010111;
        iny = 11010100;
        #100;


        inx = 10000100;
        iny = 11111110;
        #100;


        inx = 01000011;
        iny = 10101101;
        #100;


        inx = 01010100;
        iny = 00101000;
        #100;


        inx = 11010111;
        iny = 00110101;
        #100;


        inx = 01010110;
        iny = 10100100;
        #100;


        inx = 11010011;
        iny = 11101010;
        #100;


        inx = 11010101;
        iny = 00010010;
        #100;


        inx = 10001111;
        iny = 11111100;
        #100;


        inx = 11000000;
        iny = 00100110;
        #100;


        inx = 00100001;
        iny = 11110010;
        #100;


        inx = 00111100;
        iny = 10000000;
        #100;


        inx = 00111001;
        iny = 11101011;
        #100;


        inx = 11011100;
        iny = 00010100;
        #100;


        inx = 10010011;
        iny = 01011110;
        #100;


        inx = 11001110;
        iny = 10000000;
        #100;


        inx = 01111001;
        iny = 10000100;
        #100;


        inx = 01111110;
        iny = 00110100;
        #100;


        inx = 01101000;
        iny = 01001000;
        #100;


        inx = 10000111;
        iny = 00011011;
        #100;


        inx = 00100110;
        iny = 01101011;
        #100;


        inx = 01000101;
        iny = 11111110;
        #100;


        inx = 01000001;
        iny = 10101000;
        #100;


        inx = 10111110;
        iny = 10111010;
        #100;


        inx = 10111000;
        iny = 01010010;
        #100;


        inx = 10000111;
        iny = 10001011;
        #100;


        inx = 01011010;
        iny = 11111100;
        #100;


        inx = 10101111;
        iny = 00011110;
        #100;


        inx = 00110010;
        iny = 01100111;
        #100;


        inx = 10010001;
        iny = 10001011;
        #100;


        inx = 11110110;
        iny = 10111001;
        #100;


        inx = 11011110;
        iny = 10011100;
        #100;


        inx = 10111101;
        iny = 10010101;
        #100;


        inx = 00101101;
        iny = 10111001;
        #100;


        inx = 10100000;
        iny = 10101101;
        #100;


        inx = 10001010;
        iny = 00011011;
        #100;


        inx = 11101111;
        iny = 10010010;
        #100;


        inx = 11011000;
        iny = 00100111;
        #100;


        inx = 11001000;
        iny = 10010110;
        #100;


        inx = 00010100;
        iny = 10010010;
        #100;


        inx = 10011111;
        iny = 10000111;
        #100;


        inx = 00111110;
        iny = 10110001;
        #100;


        inx = 10011001;
        iny = 11001100;
        #100;


        inx = 11011000;
        iny = 11111001;
        #100;


        inx = 11011011;
        iny = 11010000;
        #100;


        inx = 00010100;
        iny = 01111100;
        #100;


        inx = 01000000;
        iny = 10011001;
        #100;


        inx = 00001010;
        iny = 11111110;
        #100;


        inx = 10010000;
        iny = 10111011;
        #100;


        inx = 11010100;
        iny = 10011111;
        #100;


        inx = 01010011;
        iny = 10010100;
        #100;


        inx = 11111100;
        iny = 11100100;
        #100;


        inx = 01001000;
        iny = 01110100;
        #100;


        inx = 11001000;
        iny = 10101000;
        #100;


        inx = 11001111;
        iny = 00100010;
        #100;


        inx = 11110000;
        iny = 00001110;
        #100;


        inx = 11110110;
        iny = 11100011;
        #100;


        inx = 11010010;
        iny = 11011100;
        #100;


        inx = 10100100;
        iny = 00000111;
        #100;


        inx = 00011010;
        iny = 11101110;
        #100;


        inx = 10010111;
        iny = 10000100;
        #100;


        inx = 01000101;
        iny = 11110010;
        #100;


        inx = 11110100;
        iny = 10000011;
        #100;


        inx = 10011110;
        iny = 11001110;
        #100;


        inx = 11111011;
        iny = 01100111;
        #100;


        inx = 10011100;
        iny = 10011010;
        #100;


        inx = 10111100;
        iny = 11110111;
        #100;


        inx = 10010100;
        iny = 10001101;
        #100;


        inx = 11001001;
        iny = 11011001;
        #100;


        inx = 11110111;
        iny = 10110001;
        #100;


        inx = 11101111;
        iny = 10010010;
        #100;


        inx = 00011001;
        iny = 11101001;
        #100;


        inx = 00011111;
        iny = 01101101;
        #100;


        inx = 00110011;
        iny = 10010000;
        #100;


        inx = 00110000;
        iny = 00001110;
        #100;


        inx = 10101110;
        iny = 11001101;
        #100;


        inx = 11001001;
        iny = 10010001;
        #100;


        inx = 01100101;
        iny = 00111101;
        #100;


        inx = 11000000;
        iny = 01000010;
        #100;


        inx = 00100101;
        iny = 01001011;
        #100;


        inx = 01100000;
        iny = 11110000;
        #100;


        inx = 01110011;
        iny = 00001101;
        #100;


        inx = 10011110;
        iny = 11011010;
        #100;


        inx = 00111001;
        iny = 01000001;
        #100;


        inx = 00101111;
        iny = 11110000;
        #100;


        inx = 11001101;
        iny = 01001101;
        #100;


        inx = 11111100;
        iny = 11011100;
        #100;


        inx = 11100011;
        iny = 00100110;
        #100;


        inx = 11000011;
        iny = 11110101;
        #100;


        inx = 11110001;
        iny = 00101000;
        #100;


        inx = 00110111;
        iny = 00001110;
        #100;


        inx = 10101000;
        iny = 10110100;
        #100;


        inx = 01110111;
        iny = 01110010;
        #100;


        inx = 11101110;
        iny = 10001011;
        #100;


        inx = 10001011;
        iny = 01110111;
        #100;


        inx = 10000001;
        iny = 01110111;
        #100;


        inx = 01101101;
        iny = 01111110;
        #100;


        inx = 11100001;
        iny = 11100000;
        #100;


        inx = 10001001;
        iny = 10001111;
        #100;


        inx = 11001100;
        iny = 11101100;
        #100;


        inx = 11011011;
        iny = 11010011;
        #100;


        inx = 11010111;
        iny = 10001110;
        #100;


        inx = 10000001;
        iny = 00000100;
        #100;


        inx = 00000000;
        iny = 01110010;
        #100;


        inx = 01110001;
        iny = 10001110;
        #100;


        inx = 11111011;
        iny = 11011100;
        #100;


        inx = 11100101;
        iny = 11110000;
        #100;


        inx = 01100110;
        iny = 01010010;
        #100;


        inx = 00101001;
        iny = 00101000;
        #100;


        inx = 11000011;
        iny = 00101110;
        #100;


        inx = 11001000;
        iny = 11101101;
        #100;


        inx = 01011000;
        iny = 01011110;
        #100;


        inx = 00100000;
        iny = 11011001;
        #100;


        inx = 11110101;
        iny = 01110001;
        #100;


        inx = 11000100;
        iny = 10101010;
        #100;


        inx = 11000111;
        iny = 01001010;
        #100;


        inx = 00111010;
        iny = 00011000;
        #100;


        inx = 01110111;
        iny = 00101111;
        #100;


        inx = 10111001;
        iny = 10100111;
        #100;


        inx = 10000100;
        iny = 11100000;
        #100;


        inx = 01011001;
        iny = 01010000;
        #100;


        inx = 10110100;
        iny = 00000001;
        #100;


        inx = 00010010;
        iny = 10001001;
        #100;


        inx = 00000001;
        iny = 11101001;
        #100;


        inx = 10011011;
        iny = 01111110;
        #100;


        inx = 00100110;
        iny = 00010111;
        #100;


        inx = 10111000;
        iny = 11001000;
        #100;


        inx = 10111101;
        iny = 01100100;
        #100;


        inx = 01101101;
        iny = 11110101;
        #100;


        inx = 01101010;
        iny = 00010101;
        #100;


        inx = 11011000;
        iny = 11100110;
        #100;


        inx = 10001100;
        iny = 00000111;
        #100;


        inx = 11111100;
        iny = 00011100;
        #100;


        inx = 11000000;
        iny = 10001101;
        #100;


        inx = 10011000;
        iny = 11111000;
        #100;


        inx = 11001011;
        iny = 00000100;
        #100;


        inx = 00001101;
        iny = 10011001;
        #100;


        inx = 00101100;
        iny = 00000010;
        #100;


        inx = 01011100;
        iny = 11000011;
        #100;


        inx = 01101010;
        iny = 10111101;
        #100;


        inx = 10010110;
        iny = 11111011;
        #100;


        inx = 00000110;
        iny = 10010110;
        #100;


        inx = 10000100;
        iny = 11011101;
        #100;


        inx = 10001010;
        iny = 01101000;
        #100;


        inx = 10100011;
        iny = 10011010;
        #100;


        inx = 10111100;
        iny = 01000000;
        #100;


        inx = 10111010;
        iny = 11101010;
        #100;


        inx = 11111101;
        iny = 10110010;
        #100;


        inx = 10001011;
        iny = 01011111;
        #100;


        inx = 11011001;
        iny = 11010100;
        #100;


        inx = 01110101;
        iny = 11100110;
        #100;


        inx = 11111111;
        iny = 10111101;
        #100;


        inx = 10001111;
        iny = 00000010;
        #100;


        inx = 10110100;
        iny = 01000011;
        #100;


        inx = 10001100;
        iny = 10011110;
        #100;


        inx = 01100110;
        iny = 10101010;
        #100;


        inx = 00011101;
        iny = 01010001;
        #100;


        inx = 11111010;
        iny = 01110110;
        #100;


        inx = 00100001;
        iny = 01000110;
        #100;


        inx = 01000000;
        iny = 00111001;
        #100;


        inx = 01100011;
        iny = 10100001;
        #100;


        inx = 10011000;
        iny = 10000111;
        #100;


        inx = 10011110;
        iny = 11101001;
        #100;


        inx = 11000011;
        iny = 11000010;
        #100;


        inx = 11001010;
        iny = 01101101;
        #100;


        inx = 01111000;
        iny = 11000001;
        #100;


        inx = 01110011;
        iny = 10001010;
        #100;


        inx = 11000101;
        iny = 10001010;
        #100;


        inx = 10111001;
        iny = 01011000;
        #100;


        inx = 10000101;
        iny = 11111111;
        #100;


        inx = 11100000;
        iny = 10101000;
        #100;


        inx = 10010010;
        iny = 11101010;
        #100;


        inx = 01111000;
        iny = 00001011;
        #100;


        inx = 10001111;
        iny = 01100001;
        #100;


        inx = 01011000;
        iny = 11000000;
        #100;


        inx = 01000011;
        iny = 10111100;
        #100;


        inx = 11011000;
        iny = 11010011;
        #100;


        inx = 11101000;
        iny = 10011111;
        #100;


        inx = 01110001;
        iny = 01011110;
        #100;


        inx = 11001100;
        iny = 00110101;
        #100;


        inx = 10000100;
        iny = 10000101;
        #100;


        inx = 10000100;
        iny = 01111110;
        #100;


        inx = 00100110;
        iny = 00111001;
        #100;


        inx = 00010100;
        iny = 11110010;
        #100;


        inx = 11001011;
        iny = 11001010;
        #100;


        inx = 01111001;
        iny = 00101000;
        #100;


        inx = 01011010;
        iny = 11100001;
        #100;


        inx = 00011000;
        iny = 11110111;
        #100;


        inx = 10101110;
        iny = 00111111;
        #100;


        inx = 01011100;
        iny = 00010101;
        #100;


        inx = 10101110;
        iny = 00111111;
        #100;


        inx = 11011110;
        iny = 01111001;
        #100;


        inx = 10000000;
        iny = 01010000;
        #100;


        inx = 10010010;
        iny = 11100100;
        #100;


        inx = 10011100;
        iny = 10000011;
        #100;


        inx = 01101110;
        iny = 01000010;
        #100;


        inx = 10010100;
        iny = 00001111;
        #100;


        inx = 10111101;
        iny = 00111111;
        #100;


        inx = 10100110;
        iny = 10010111;
        #100;


        inx = 01011101;
        iny = 01001111;
        #100;


        inx = 01110010;
        iny = 10010011;
        #100;


        inx = 00111111;
        iny = 11010101;
        #100;


        inx = 10001010;
        iny = 01000110;
        #100;


        inx = 10001001;
        iny = 00001101;
        #100;


        inx = 10000011;
        iny = 11110000;
        #100;


        inx = 11111011;
        iny = 00000110;
        #100;


        inx = 00110010;
        iny = 00101101;
        #100;


        inx = 10000000;
        iny = 01111110;
        #100;


        inx = 11101111;
        iny = 00100100;
        #100;


        inx = 00111011;
        iny = 11101011;
        #100;


        inx = 00111010;
        iny = 11110100;
        #100;


        inx = 01100100;
        iny = 00100100;
        #100;


        inx = 11010010;
        iny = 01110001;
        #100;


        inx = 00100001;
        iny = 01110001;
        #100;


        inx = 01111010;
        iny = 00000111;
        #100;


        inx = 00111010;
        iny = 00010100;
        #100;


        inx = 10001101;
        iny = 00101111;
        #100;


        inx = 00000000;
        iny = 11101010;
        #100;


        inx = 11110100;
        iny = 01000100;
        #100;


        inx = 00001000;
        iny = 01011101;
        #100;


        inx = 10111110;
        iny = 10101110;
        #100;


        inx = 11000111;
        iny = 10000011;
        #100;


        inx = 10000111;
        iny = 11110111;
        #100;


        inx = 10111001;
        iny = 01111111;
        #100;


        inx = 10101000;
        iny = 10111111;
        #100;


        inx = 01001011;
        iny = 11011110;
        #100;


        inx = 00100110;
        iny = 00000111;
        #100;


        inx = 01010111;
        iny = 10001100;
        #100;


        inx = 10001000;
        iny = 01101100;
        #100;


        inx = 11011110;
        iny = 01101110;
        #100;


        inx = 10111011;
        iny = 11111001;
        #100;


        inx = 00011011;
        iny = 11110010;
        #100;


        inx = 11000000;
        iny = 00111111;
        #100;


        inx = 11111100;
        iny = 01001000;
        #100;


        inx = 01110101;
        iny = 11000111;
        #100;


        inx = 10001011;
        iny = 10111100;
        #100;


        inx = 10111001;
        iny = 11111110;
        #100;


        inx = 10101100;
        iny = 11110100;
        #100;


        inx = 11111001;
        iny = 11100011;
        #100;


        inx = 00111111;
        iny = 10011000;
        #100;


        inx = 01001100;
        iny = 11111111;
        #100;


        inx = 01111010;
        iny = 00001010;
        #100;


        inx = 10110010;
        iny = 01101011;
        #100;


        inx = 01111110;
        iny = 01111011;
        #100;


        inx = 01011101;
        iny = 00011001;
        #100;


        inx = 11000101;
        iny = 00101010;
        #100;


        inx = 11100111;
        iny = 01111010;
        #100;


        inx = 11011001;
        iny = 10100101;
        #100;


        inx = 00001111;
        iny = 10110000;
        #100;


        inx = 10110000;
        iny = 00000111;
        #100;


        inx = 10010001;
        iny = 01000000;
        #100;


        inx = 11101011;
        iny = 10101101;
        #100;


        inx = 01100001;
        iny = 11001101;
        #100;


        inx = 01000011;
        iny = 01111010;
        #100;


        inx = 00001100;
        iny = 10001101;
        #100;


        inx = 00010000;
        iny = 01000110;
        #100;


        inx = 11110111;
        iny = 00100100;
        #100;


        inx = 11011111;
        iny = 01011110;
        #100;


        inx = 00011001;
        iny = 11100000;
        #100;


        inx = 10110111;
        iny = 11110100;
        #100;


        inx = 00001110;
        iny = 10001001;
        #100;


        inx = 00110001;
        iny = 10001010;
        #100;


        inx = 11111111;
        iny = 10111110;
        #100;


        inx = 01110000;
        iny = 00000100;
        #100;


        inx = 10110110;
        iny = 11100100;
        #100;


        inx = 11000001;
        iny = 01111000;
        #100;


        inx = 10011011;
        iny = 01111100;
        #100;


        inx = 01101010;
        iny = 01100111;
        #100;


        inx = 00010100;
        iny = 11011000;
        #100;


        inx = 01011010;
        iny = 10100110;
        #100;


        inx = 00111000;
        iny = 01111111;
        #100;


        inx = 10011010;
        iny = 01100101;
        #100;


        inx = 11001011;
        iny = 00001001;
        #100;


        inx = 00010111;
        iny = 11110011;
        #100;


        inx = 10100000;
        iny = 01110110;
        #100;


        inx = 00011111;
        iny = 11010100;
        #100;


        inx = 10100011;
        iny = 10010110;
        #100;


        inx = 10000010;
        iny = 11001111;
        #100;


        inx = 11011010;
        iny = 11101010;
        #100;


        inx = 11011001;
        iny = 10111111;
        #100;


        inx = 00011110;
        iny = 01110101;
        #100;


        inx = 10011001;
        iny = 00000111;
        #100;


        inx = 00111110;
        iny = 10100010;
        #100;


        inx = 10111011;
        iny = 10100001;
        #100;


        inx = 11110000;
        iny = 10011011;
        #100;


        inx = 11101110;
        iny = 01000100;
        #100;


        inx = 10111010;
        iny = 00110011;
        #100;


        inx = 10101010;
        iny = 01010100;
        #100;


        inx = 01001001;
        iny = 00011011;
        #100;


        inx = 11001111;
        iny = 10001001;
        #100;


        inx = 10010111;
        iny = 10000110;
        #100;


        inx = 00001101;
        iny = 01011000;
        #100;


        inx = 00111011;
        iny = 11011101;
        #100;


        inx = 00010001;
        iny = 10011111;
        #100;


        inx = 01111111;
        iny = 01110110;
        #100;


        inx = 00110111;
        iny = 10000010;
        #100;


        inx = 00010011;
        iny = 10010101;
        #100;


        inx = 11100101;
        iny = 00011110;
        #100;


        inx = 11010111;
        iny = 01011110;
        #100;


        inx = 00111110;
        iny = 01011110;
        #100;


        inx = 11001110;
        iny = 10100111;
        #100;


        inx = 01111111;
        iny = 11101100;
        #100;


        inx = 10010100;
        iny = 01111010;
        #100;


        inx = 11110110;
        iny = 01100100;
        #100;


        inx = 01000100;
        iny = 00001111;
        #100;


        inx = 10100110;
        iny = 01010110;
        #100;


        inx = 10111110;
        iny = 01110101;
        #100;


        inx = 01110111;
        iny = 11101111;
        #100;


        inx = 01010110;
        iny = 01001011;
        #100;


        inx = 00101011;
        iny = 01101011;
        #100;


        inx = 10001001;
        iny = 11110000;
        #100;


        inx = 11010011;
        iny = 00010111;
        #100;


        inx = 01001101;
        iny = 10000011;
        #100;


        inx = 00110000;
        iny = 00000011;
        #100;


        inx = 00100110;
        iny = 11001011;
        #100;


        inx = 11111110;
        iny = 01101110;
        #100;


        inx = 11011111;
        iny = 00011110;
        #100;


        inx = 00111100;
        iny = 01100001;
        #100;


        inx = 11111010;
        iny = 01100001;
        #100;


        inx = 10000101;
        iny = 10000110;
        #100;


        inx = 01101100;
        iny = 00001100;
        #100;


        inx = 01011011;
        iny = 01101000;
        #100;


        inx = 10001110;
        iny = 01010010;
        #100;


        inx = 00110111;
        iny = 10001101;
        #100;


        inx = 11001010;
        iny = 00100011;
        #100;


        inx = 11111111;
        iny = 11101001;
        #100;


        inx = 00101001;
        iny = 10010001;
        #100;


        inx = 01001110;
        iny = 11000000;
        #100;


        inx = 01101110;
        iny = 11010110;
        #100;


        inx = 00000110;
        iny = 01010111;
        #100;


        inx = 10001110;
        iny = 10110111;
        #100;


        inx = 00101111;
        iny = 11000100;
        #100;


        inx = 00101100;
        iny = 00111110;
        #100;


        inx = 10011011;
        iny = 01100010;
        #100;


        inx = 10001010;
        iny = 00101011;
        #100;


        inx = 00001101;
        iny = 01100101;
        #100;


        inx = 00110010;
        iny = 01111010;
        #100;


        inx = 01100111;
        iny = 00111000;
        #100;


        inx = 10110001;
        iny = 10001111;
        #100;


        inx = 11010011;
        iny = 10100110;
        #100;


        inx = 10110010;
        iny = 00100101;
        #100;


        inx = 10111111;
        iny = 00010001;
        #100;


        inx = 00011011;
        iny = 10110010;
        #100;


        inx = 10011010;
        iny = 11001111;
        #100;


        inx = 01101000;
        iny = 00010111;
        #100;


        inx = 10011011;
        iny = 11111000;
        #100;


        inx = 11001001;
        iny = 10010110;
        #100;


        inx = 01011110;
        iny = 10010110;
        #100;


        inx = 00000100;
        iny = 11001011;
        #100;


        inx = 00101100;
        iny = 11100101;
        #100;


        inx = 00000000;
        iny = 00110000;
        #100;


        inx = 00100000;
        iny = 11011110;
        #100;


        inx = 10100101;
        iny = 01100000;
        #100;


        inx = 11101010;
        iny = 00110001;
        #100;


        inx = 01110010;
        iny = 01001111;
        #100;


        inx = 01010000;
        iny = 00101010;
        #100;


        inx = 10000100;
        iny = 10101101;
        #100;


        inx = 00110000;
        iny = 00001000;
        #100;


        inx = 00111101;
        iny = 11100101;
        #100;


        inx = 11011110;
        iny = 00100101;
        #100;


        inx = 11111111;
        iny = 10011000;
        #100;


        inx = 00000111;
        iny = 01111111;
        #100;


        inx = 10111001;
        iny = 11111010;
        #100;


        inx = 10101111;
        iny = 01000110;
        #100;


        inx = 10111001;
        iny = 01001001;
        #100;


        inx = 10001001;
        iny = 10011010;
        #100;


        inx = 10101100;
        iny = 00000011;
        #100;


        inx = 00000010;
        iny = 11111011;
        #100;


        inx = 11010000;
        iny = 01100111;
        #100;


        inx = 01110001;
        iny = 00110110;
        #100;


        inx = 01001101;
        iny = 11000111;
        #100;


        inx = 11110001;
        iny = 11111100;
        #100;


        inx = 11000100;
        iny = 01110010;
        #100;


        inx = 10110010;
        iny = 10000000;
        #100;


        inx = 11111011;
        iny = 10001111;
        #100;


        inx = 10111110;
        iny = 01000110;
        #100;


        inx = 11011100;
        iny = 10001010;
        #100;


        inx = 00100111;
        iny = 00010111;
        #100;


        inx = 11011101;
        iny = 10010100;
        #100;


        inx = 11001100;
        iny = 11000010;
        #100;


        inx = 11111000;
        iny = 11111100;
        #100;


        inx = 00000110;
        iny = 10110000;
        #100;


        inx = 11001010;
        iny = 11001111;
        #100;


        inx = 11101111;
        iny = 11110011;
        #100;


        inx = 00001001;
        iny = 01000010;
        #100;


        inx = 11010011;
        iny = 01011001;
        #100;


        inx = 00100001;
        iny = 00111101;
        #100;


        inx = 00011111;
        iny = 00000001;
        #100;


        inx = 11100010;
        iny = 10110101;
        #100;


        inx = 10110111;
        iny = 01111011;
        #100;


        inx = 11101101;
        iny = 00100010;
        #100;


        inx = 00101010;
        iny = 10001110;
        #100;


        inx = 01100100;
        iny = 01100001;
        #100;


        inx = 10110010;
        iny = 10001110;
        #100;


        inx = 01101001;
        iny = 00100011;
        #100;


        inx = 00110100;
        iny = 11011011;
        #100;


        inx = 11010011;
        iny = 01010010;
        #100;


        inx = 10110111;
        iny = 11000110;
        #100;


        inx = 00011001;
        iny = 10010010;
        #100;


        inx = 01110000;
        iny = 01110110;
        #100;


        inx = 10111000;
        iny = 10111110;
        #100;


        inx = 10001111;
        iny = 11101110;
        #100;


        inx = 01010010;
        iny = 01000010;
        #100;


        inx = 01001110;
        iny = 11101101;
        #100;


        inx = 10000010;
        iny = 11010100;
        #100;


        inx = 11010001;
        iny = 00001101;
        #100;


        inx = 10000111;
        iny = 00111000;
        #100;


        inx = 01100000;
        iny = 11101100;
        #100;


        inx = 11111010;
        iny = 01101111;
        #100;


        inx = 01101001;
        iny = 11101001;
        #100;


        inx = 00001000;
        iny = 10100011;
        #100;


        inx = 00001000;
        iny = 01001110;
        #100;


        inx = 00001111;
        iny = 11101101;
        #100;


        inx = 00110110;
        iny = 10011100;
        #100;


        inx = 01110000;
        iny = 10011100;
        #100;


        inx = 10100011;
        iny = 10101100;
        #100;


        inx = 00101001;
        iny = 11100100;
        #100;


        inx = 11011110;
        iny = 00100100;
        #100;


        inx = 10010010;
        iny = 01010011;
        #100;


        inx = 10101011;
        iny = 11111110;
        #100;


        inx = 00011010;
        iny = 00011111;
        #100;


        inx = 11010110;
        iny = 01101000;
        #100;


        inx = 01101110;
        iny = 11101011;
        #100;


        inx = 01000111;
        iny = 10001011;
        #100;


        inx = 11101110;
        iny = 10010010;
        #100;


        inx = 00011000;
        iny = 00111111;
        #100;


        inx = 11001101;
        iny = 10011001;
        #100;


        inx = 00100101;
        iny = 01100101;
        #100;


        inx = 11110110;
        iny = 10010001;
        #100;


        inx = 01111100;
        iny = 00001011;
        #100;


        inx = 00010111;
        iny = 10110100;
        #100;


        inx = 00111000;
        iny = 10111000;
        #100;


        inx = 01000011;
        iny = 11111101;
        #100;


        inx = 11011110;
        iny = 00111100;
        #100;


        inx = 00111101;
        iny = 11001001;
        #100;


        inx = 10101011;
        iny = 11101111;
        #100;


        inx = 11101010;
        iny = 10000001;
        #100;


        inx = 00001000;
        iny = 01110000;
        #100;


        inx = 01001101;
        iny = 11010101;
        #100;


        inx = 11101101;
        iny = 10100011;
        #100;


        inx = 10010001;
        iny = 10100011;
        #100;


        inx = 11110101;
        iny = 10001001;
        #100;


        inx = 11001001;
        iny = 10101110;
        #100;


        inx = 10000100;
        iny = 00101111;
        #100;


        inx = 00000101;
        iny = 10100001;
        #100;


        inx = 00001100;
        iny = 01110011;
        #100;


        inx = 10001101;
        iny = 11111011;
        #100;


        inx = 10010010;
        iny = 00101001;
        #100;


        inx = 11111110;
        iny = 01110111;
        #100;


        inx = 10110111;
        iny = 10111000;
        #100;


        inx = 01111000;
        iny = 00001001;
        #100;


        inx = 01100111;
        iny = 11001100;
        #100;


        inx = 10100110;
        iny = 10101011;
        #100;


        inx = 01000101;
        iny = 01101000;
        #100;


        inx = 11011000;
        iny = 00010001;
        #100;


        inx = 01110011;
        iny = 00100010;
        #100;


        inx = 01100100;
        iny = 00011110;
        #100;


        inx = 11101101;
        iny = 01100011;
        #100;


        inx = 11010110;
        iny = 00101100;
        #100;


        inx = 10000011;
        iny = 10110111;
        #100;


        inx = 01001010;
        iny = 11110100;
        #100;


        inx = 00111101;
        iny = 00101100;
        #100;


        inx = 01001011;
        iny = 01000110;
        #100;


        inx = 11110111;
        iny = 10011001;
        #100;


        inx = 00011011;
        iny = 00001101;
        #100;


        inx = 11111110;
        iny = 01000110;
        #100;


        inx = 00010110;
        iny = 01100101;
        #100;


        inx = 01101110;
        iny = 01110001;
        #100;


        inx = 00100010;
        iny = 11101000;
        #100;


        inx = 00100111;
        iny = 10000100;
        #100;


        inx = 01111110;
        iny = 00011000;
        #100;


        inx = 01001000;
        iny = 00001101;
        #100;


        inx = 01111111;
        iny = 01100010;
        #100;


        inx = 01010001;
        iny = 00000111;
        #100;


        inx = 00101010;
        iny = 01100110;
        #100;


        inx = 10000110;
        iny = 01010111;
        #100;


        inx = 00000010;
        iny = 01010100;
        #100;


        inx = 11100110;
        iny = 00010011;
        #100;


        inx = 00011111;
        iny = 11100000;
        #100;


        inx = 01110111;
        iny = 11000111;
        #100;


        inx = 10001100;
        iny = 11111010;
        #100;


        inx = 10110101;
        iny = 10011101;
        #100;


        inx = 10111110;
        iny = 10010101;
        #100;


        inx = 00000001;
        iny = 00110110;
        #100;


        inx = 01000110;
        iny = 00000101;
        #100;


        inx = 10101111;
        iny = 10001001;
        #100;


        inx = 11000000;
        iny = 01001101;
        #100;


        inx = 10111000;
        iny = 00110010;
        #100;


        inx = 01010001;
        iny = 00000000;
        #100;


        inx = 00100011;
        iny = 00000011;
        #100;


        inx = 00111000;
        iny = 00001101;
        #100;


        inx = 01001100;
        iny = 11011011;
        #100;


        inx = 00000101;
        iny = 10011100;
        #100;


        inx = 11111000;
        iny = 00010010;
        #100;


        inx = 00100001;
        iny = 00011110;
        #100;


        inx = 01000101;
        iny = 10000111;
        #100;


        inx = 01101101;
        iny = 10001111;
        #100;


        inx = 00001011;
        iny = 00101101;
        #100;


        inx = 11101110;
        iny = 10010000;
        #100;


        inx = 00011100;
        iny = 01000101;
        #100;


        inx = 01001100;
        iny = 10001110;
        #100;


        inx = 10001001;
        iny = 11100100;
        #100;


        inx = 10101001;
        iny = 01100000;
        #100;


        inx = 10100101;
        iny = 00100110;
        #100;


        inx = 01100010;
        iny = 11110000;
        #100;


        inx = 00001001;
        iny = 10010011;
        #100;


        inx = 11110010;
        iny = 01101011;
        #100;


        inx = 00110111;
        iny = 11110110;
        #100;


        inx = 00111000;
        iny = 10000000;
        #100;


        inx = 01101110;
        iny = 11001000;
        #100;


        inx = 10101011;
        iny = 00001110;
        #100;


        inx = 01111000;
        iny = 01011110;
        #100;


        inx = 00100010;
        iny = 01001000;
        #100;


        inx = 01011010;
        iny = 00101001;
        #100;


        inx = 10111011;
        iny = 10011101;
        #100;


        inx = 01100010;
        iny = 10101001;
        #100;


        inx = 01111000;
        iny = 10000001;
        #100;


        inx = 00001110;
        iny = 01001101;
        #100;


        inx = 11011111;
        iny = 00111000;
        #100;


        inx = 00010010;
        iny = 00011010;
        #100;


        inx = 10111110;
        iny = 11001111;
        #100;


        inx = 01011010;
        iny = 00101110;
        #100;


        inx = 01011101;
        iny = 01101110;
        #100;


        inx = 00011011;
        iny = 11010001;
        #100;


        inx = 10001011;
        iny = 01001101;
        #100;


        inx = 11011011;
        iny = 00111011;
        #100;


        inx = 01111010;
        iny = 10100011;
        #100;


        inx = 10010010;
        iny = 00001010;
        #100;


        inx = 10011001;
        iny = 11101010;
        #100;


        inx = 10100110;
        iny = 01110101;
        #100;


        inx = 01111010;
        iny = 00111111;
        #100;


        inx = 11110001;
        iny = 01010011;
        #100;


        inx = 10011011;
        iny = 01010101;
        #100;


        inx = 10101011;
        iny = 10010001;
        #100;


        inx = 10000000;
        iny = 10010011;
        #100;


        inx = 11111101;
        iny = 10011011;
        #100;


        inx = 10001101;
        iny = 10101001;
        #100;


        inx = 00110010;
        iny = 10001011;
        #100;


        inx = 11001010;
        iny = 11100001;
        #100;


        inx = 01000001;
        iny = 11111111;
        #100;


        inx = 11011001;
        iny = 01010001;
        #100;


        inx = 01111000;
        iny = 00110010;
        #100;


        inx = 01111110;
        iny = 11011001;
        #100;


        inx = 00100110;
        iny = 10100100;
        #100;


        inx = 00000101;
        iny = 00011011;
        #100;


        inx = 00100101;
        iny = 10100111;
        #100;


        inx = 11110001;
        iny = 01111010;
        #100;


        inx = 00000000;
        iny = 01111011;
        #100;


        inx = 00010011;
        iny = 10100111;
        #100;


        inx = 10101100;
        iny = 00101000;
        #100;


        inx = 00001110;
        iny = 10011110;
        #100;


        inx = 11010111;
        iny = 10100010;
        #100;


        inx = 11011011;
        iny = 00011000;
        #100;


        inx = 00111000;
        iny = 11101101;
        #100;


        inx = 00101010;
        iny = 01001111;
        #100;


        inx = 01100010;
        iny = 01011010;
        #100;


        inx = 01110100;
        iny = 10110101;
        #100;


        inx = 11111111;
        iny = 00010000;
        #100;


        inx = 11110011;
        iny = 11100110;
        #100;


        inx = 11001000;
        iny = 00010001;
        #100;


        inx = 11111110;
        iny = 00010010;
        #100;


        inx = 01100001;
        iny = 10000100;
        #100;


        inx = 00101000;
        iny = 00110101;
        #100;


        inx = 11101100;
        iny = 10110010;
        #100;


        inx = 00010001;
        iny = 11101101;
        #100;


        inx = 01110101;
        iny = 01010100;
        #100;


        inx = 10000111;
        iny = 01100000;
        #100;


        inx = 01101101;
        iny = 10000000;
        #100;


        inx = 11001010;
        iny = 10111000;
        #100;


        inx = 11100011;
        iny = 00110100;
        #100;


        inx = 01100000;
        iny = 00000010;
        #100;


        inx = 00100000;
        iny = 11101000;
        #100;


        inx = 00000001;
        iny = 01000111;
        #100;


        inx = 10101001;
        iny = 10011000;
        #100;


        inx = 01011101;
        iny = 11000101;
        #100;


        inx = 01010000;
        iny = 11001110;
        #100;


        inx = 10100110;
        iny = 11110111;
        #100;


        inx = 11110111;
        iny = 10101000;
        #100;


        inx = 00111110;
        iny = 01111111;
        #100;


        inx = 01011100;
        iny = 11110010;
        #100;


        inx = 11110001;
        iny = 11000011;
        #100;


        inx = 00111001;
        iny = 00000111;
        #100;


        inx = 00000011;
        iny = 10100110;
        #100;


        inx = 11000001;
        iny = 10110011;
        #100;


        inx = 10000000;
        iny = 10100111;
        #100;


        inx = 10000011;
        iny = 01100000;
        #100;


        inx = 00010111;
        iny = 01000111;
        #100;


        inx = 11000010;
        iny = 01100110;
        #100;


        inx = 11111110;
        iny = 00101110;
        #100;


        inx = 11001011;
        iny = 00000111;
        #100;


        inx = 11011010;
        iny = 10110000;
        #100;


        inx = 01001001;
        iny = 10100101;
        #100;


        inx = 10110001;
        iny = 00110101;
        #100;


        inx = 10110100;
        iny = 01010110;
        #100;


        inx = 11111101;
        iny = 00110011;
        #100;


        inx = 01111101;
        iny = 01111110;
        #100;


        inx = 10000101;
        iny = 10101000;
        #100;


        inx = 00100011;
        iny = 11101001;
        #100;


        inx = 01001010;
        iny = 11010011;
        #100;


        inx = 01010111;
        iny = 00101110;
        #100;


        inx = 10010111;
        iny = 01111100;
        #100;


        inx = 00101011;
        iny = 10001010;
        #100;


        inx = 11111010;
        iny = 10001111;
        #100;


        inx = 11100010;
        iny = 00101100;
        #100;


        inx = 11010011;
        iny = 10011011;
        #100;


        inx = 01110010;
        iny = 01111101;
        #100;


        inx = 10110100;
        iny = 00010110;
        #100;


        inx = 10010011;
        iny = 01010001;
        #100;


        inx = 00110101;
        iny = 01111011;
        #100;


        inx = 10101000;
        iny = 11111000;
        #100;


        inx = 01100100;
        iny = 00000000;
        #100;


        inx = 11000101;
        iny = 10000111;
        #100;


        inx = 10110000;
        iny = 00111000;
        #100;


        inx = 11101111;
        iny = 11110011;
        #100;


        inx = 10100010;
        iny = 00101111;
        #100;


        inx = 01110001;
        iny = 00011011;
        #100;


        inx = 01111101;
        iny = 10011101;
        #100;


        inx = 00100011;
        iny = 00001100;
        #100;


    end
endmodule
